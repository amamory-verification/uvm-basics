interface dut_if();

	logic clock, reset;
	logic dout;
endinterface : dut_if
