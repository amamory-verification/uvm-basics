class hermes_noc_seq_config extends uvm_object;
`uvm_object_utils(hermes_noc_seq_config)


//==========================
// seq item knobs
//==========================
// set the input router port where the sequence will inject its packets. default is 0  
//rand bit [4:0] source_router;
// set the random distribution for port 
bit [4:0] router_dist[hermes_pkg::NROT] = {1,1,1,1,1,1,1,1,1};

/*
constraint c_router {
  source_router inside { [0:hermes_pkg::NROT-1] };
  source_router dist { 
  	0 := router_dist[0],
  	1 := router_dist[1],
  	2 := router_dist[2],
  	3 := router_dist[3],
  	4 := router_dist[4],
    5 := router_dist[5],
    6 := router_dist[6],
    7 := router_dist[7],
    8 := router_dist[8]
  };
}
*/

// set the packet size
rand hermes_packet_t::packet_size_t p_size;
// weights for packet size
bit [4:0] w_zero=1, w_small=2, w_med=10, w_large=1;

// choose random packet size with weights
constraint c_p_size {
  p_size dist {
    //hermes_packet_t::ZERO  := w_zero, // not supported by the router. enable only to generated invalid packets
    hermes_packet_t::SMALL := w_small,
    hermes_packet_t::MED   := w_med,
    hermes_packet_t::LARGE := w_large
  };
}

// target packet address
rand bit [7:0] header;

constraint c_header { 
  // the possible target address
  header inside {8'h00,8'h01,8'h02,8'h10, 8'h11,8'h12,8'h20, 8'h21,8'h22};
}

//==========================
// seq knobs 
//==========================
// set the # of packets generated by the sequence
rand int npackets = 1;

constraint c_packets { 
  npackets inside {[1:200]};
  npackets dist   { 
      [1:20]    := 20, 
      [21:50]   := 10, 
      [51:100]  := 5, 
      [101:200] := 1
  };
}


function void do_copy( uvm_object rhs );
  hermes_noc_seq_config that;

  if ( ! $cast( that, rhs ) ) begin
     `uvm_error( get_name(), "rhs is not a hermes_noc_seq_config" )
     return;
  end

  super.do_copy( rhs );
  //this.source_router   = that.source_router;
  this.router_dist     = that.router_dist;
  this.p_size          = that.p_size;
  this.w_zero          = that.w_zero;
  this.w_small         = that.w_small;
  this.w_med           = that.w_med;
  this.w_large         = that.w_large;
  this.header          = that.header;
  this.npackets        = that.npackets;
endfunction: do_copy


virtual function string convert2string();
  string s = super.convert2string();      
  //s = { s, $psprintf( "\n port       : %0d", source_router) };
  s = { s, $psprintf( "\n p_size     : %0d", p_size) };
  s = { s, $psprintf( "\n header     : %H" , header) };
  //s = { s, $psprintf( "\n valid_addr : %p" , hermes_pkg::valid_addrs(port)) };
  s = { s, $psprintf( "\n npackets   : %0d", npackets) };
  return s;
endfunction: convert2string

function new( string name = "" );
  super.new( name );
endfunction: new

endclass
