package my_sequences;


class seq_of_commands extends uvm_sequence #(my_transaction);

class read_modify_write extends uvm_sequence #(my_transaction);

class my_sequence extends uvm_sequence #(my_transaction);


endpackage
