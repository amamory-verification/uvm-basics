/*
 this flat sequence injects 'npackets' into a single port 'port'   
*/
class basic_seq extends base_vseq; 
`uvm_object_utils(basic_seq)


function new(string name = "basic_seq");
  super.new(name);
endfunction: new

//==========================
// seq item knobs
//==========================
rand packet_t::packet_size_t p_size;
// weights for packet size
bit [4:0] w_zero=1, w_small=2, w_med=10, w_large=1;

// choose random packet size with weights
constraint c_p_size {
  p_size dist {
    packet_t::ZERO  := w_zero,
    packet_t::SMALL := w_small,
    packet_t::MED   := w_med,
    packet_t::LARGE := w_large
  };
}


// target packet address
rand bit [7:0] header;
// it contains the valid target addresses
bit [7:0] valid_target_addr[$];

constraint c_header { 
  header inside {valid_target_addr};
}

//==========================
// seq item timing knobs
//==========================
// randomize the number of cycles the driver waits to start sending the packet. used by driver
rand bit [3:0] cycle2send;
// used to change the random distribution of  cycle2send
bit [3:0] cycle2send_dist[16] = {10,10,10,1,1,1,1,1,1,1,1,1,1,1,1,1};


// randomize the number of cycles between flits. used by driver
rand bit [3:0] cycle2flit;
// used to change the random distribution of  cycle2flit
bit [3:0] cycle2flit_dist[16] = {15,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1};

//==========================
// seq knobs 
//==========================
// set the # of packets generated by the sequence. default is 50
rand int npackets;

constraint c_packets { 
  npackets inside {[1:200]};
  npackets dist   { 
      [1:20]    := 20, 
      [21:50]   := 10, 
      [51:100]  := 5, 
      [101:200] := 1
  };
}


function void pre_randomize();
  valid_target_addr = router_pkg::valid_addrs(this.port);
endfunction

task body;
  packet_t tx;
  repeat(this.npackets)
  begin
    tx = packet_t::type_id::create("tx");
    // set the driver port where these packets will be injected
    tx.dport = this.port;
    // disable packets with zero payload
    tx.w_zero = 0;
    assert(tx.randomize() with {
        tx.p_size == this.p_size;
        tx.header == this.header;
        tx.cycle2send == this.cycle2send;
        tx.cycle2flit == this.cycle2flit;
      }
    );
    start_item(tx);
    // this.header is the default value, then it means that it must be randomized, else, it must use the assinged value
    /*
    if (this.header == 8'hFF) 
      assert(tx.randomize() with {tx.p_size == psize;});
    else begin
      //tx.header.mode(0);
      assert(tx.randomize() with {tx.p_size == psize; tx.header == header;});
    end
*/
    
    //assert(tx.randomize());
    //assert(tx.randomize() with {tx.payload.size() == 1;});
    finish_item(tx);
  end
endtask: body

endclass: basic_seq

