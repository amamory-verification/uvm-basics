class seq_config extends uvm_object;
`uvm_object_utils(seq_config)




//==========================
// seq item knobs
//==========================
// set the input router port where the sequence will inject its packets. default is 0  
rand bit [3:0] port;
// set the random distribution for port 
bit [3:0] port_dist[router_pkg::NPORT] = {1,1,1,1,1};

constraint c_port {
  port inside { [0:router_pkg::NPORT-1] };
  port dist { 
  	0 := port_dist[0],
  	1 := port_dist[1],
  	2 := port_dist[2],
  	3 := port_dist[3],
  	4 := port_dist[4]
  };
}

// set the packet size
rand packet_t::packet_size_t p_size;
// weights for packet size
bit [4:0] w_zero=1, w_small=2, w_med=10, w_large=1;

// choose random packet size with weights
constraint c_p_size {
  p_size dist {
    //packet_t::ZERO  := w_zero, // not supported by the router. enable only to generated invalid packets
    packet_t::SMALL := w_small,
    packet_t::MED   := w_med,
    packet_t::LARGE := w_large
  };
}


// target packet address
rand bit [7:0] header;

constraint c_header { 
  // given the input port 'port', it returns the list of possible target address for the header
  header inside {router_pkg::valid_addrs(this.port)};
  // the list of valid address depends on the input port
  solve port before header;
}


/*
//==========================
// seq item timing knobs
//==========================
// randomize the number of cycles the driver waits to start sending the packet. used by driver
rand bit [3:0] cycle2send;
// used to change the random distribution of  cycle2send
bit [3:0] cycle2send_dist[16] = {10,10,10,1,1,1,1,1,1,1,1,1,1,1,1,1};


// randomize the number of cycles between flits. used by driver
rand bit [3:0] cycle2flit;
// used to change the random distribution of  cycle2flit
bit [3:0] cycle2flit_dist[16] = {15,5,5,1,1,1,1,1,1,1,1,1,1,1,1,1};
*/

//==========================
// seq knobs 
//==========================
// set the # of packets generated by the sequence
rand int npackets = 1;

constraint c_packets { 
  npackets inside {[1:200]};
  npackets dist   { 
      [1:20]    := 20, 
      [21:50]   := 10, 
      [51:100]  := 5, 
      [101:200] := 1
  };
}


function void do_copy( uvm_object rhs );
  seq_config that;

  if ( ! $cast( that, rhs ) ) begin
     `uvm_error( get_name(), "rhs is not a seq_config" )
     return;
  end

  super.do_copy( rhs );
  this.port            = that.port;
  this.port_dist       = that.port_dist;
  this.p_size          = that.p_size;
  this.w_zero          = that.w_zero;
  this.w_small         = that.w_small;
  this.w_med           = that.w_med;
  this.w_large         = that.w_large;
  this.header          = that.header;
  //this.cycle2send      = that.cycle2send;
  //this.cycle2send_dist = that.cycle2send_dist;
  //this.cycle2flit      = that.cycle2flit;
  //this.cycle2flit_dist = that.cycle2flit_dist;
  this.npackets        = that.npackets;
endfunction: do_copy


virtual function string convert2string();
  string s = super.convert2string();      
  s = { s, $psprintf( "\n port       : %0d", port) };
  s = { s, $psprintf( "\n p_size     : %0d", p_size) };
  s = { s, $psprintf( "\n header     : %H" , header) };
  s = { s, $psprintf( "\n valid_addr : %p" , router_pkg::valid_addrs(port)) };
  //s = { s, $psprintf( "\n cycle2send : %0d", cycle2send) };
  //s = { s, $psprintf( "\n cycle2flit : %0d", cycle2flit) };
  s = { s, $psprintf( "\n npackets   : %0d", npackets) };
  return s;
endfunction: convert2string

endclass
