interface hermes_monitor_bfm(hermes_if bus);
	// TO Be DONE
endinterface