package hermes_noc_seq_pkg;

   import uvm_pkg::*;
   import hermes_pkg::*;
  
   `include "uvm_macros.svh"

   `include "src/hermes_noc_base_seq.sv"
   `include "src/hermes_noc_seq_config.sv"
   `include "src/repeat_seq.sv"
/*
   `include "src/parallel_seq.sv"
*/
endpackage
