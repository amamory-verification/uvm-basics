interface hermes_driver_bfm(hermes_if bus);
	// TO Be DONE
endinterface