----------------------------------------------------------------
--                                   CROSSBAR
--                                    --------------
--              DATA_AV ->|                 |
--              DATA_IN ->|                 |
--            DATA_ACK <-|                 |-> TX
--                 SENDER ->|                 |-> DATA_OUT
--                       FREE ->|                  |<- CREDIT_I
--                 TAB_IN ->|                  |
--              TAB_OUT ->|                  |
--                                    --------------
----------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use work.HermesPackage.all;

entity Hermes_crossbar_TC is
port(
	data_av:     in  regNport;
	data_in:     in  arrayNport_regflit;
	data_ack:    out regNport;
	sender:      in  regNport;
	free:        in  regNport;
	tab_in:      in  arrayNport_reg3;
	tab_out:     in  arrayNport_reg3;
	tx:          out regNport;
	data_out:    out arrayNport_regflit;
	credit_i:    in  regNport);
end Hermes_crossbar_TC;

architecture AlgorithmXY of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else 			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else
			 data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else 			
			credit_i(SOUTH) when tab_in(WEST)="011" and data_av(WEST)='1' else
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';

----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_av(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_in(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmXY;
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
architecture AlgorithmWFNM of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_av(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_in(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else
			data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else			
			credit_i(SOUTH) when tab_in(WEST)="011" and data_av(WEST)='1' else
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_av(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_in(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(EAST) when tab_in(SOUTH)="000" and data_av(SOUTH)='1' else			
			credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmWFNM;
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
architecture AlgorithmNLNM of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else		
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else					
			credit_i(SOUTH) when tab_in(WEST)="011" and data_av(WEST)='1' else
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_av(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_in(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmNLNM;
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
architecture AlgorithmNFNM of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';	
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_av(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_in(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else			
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else			
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(EAST) when tab_in(SOUTH)="000" and data_av(SOUTH)='1' else			
			credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmNFNM;
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
architecture AlgorithmWFM of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_av(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_in(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else
			data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else			
			credit_i(SOUTH) when tab_in(WEST)="011" and data_av(WEST)='1' else
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_av(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_in(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(EAST) when tab_in(SOUTH)="000" and data_av(SOUTH)='1' else			
			credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmWFM;
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
architecture AlgorithmNLM of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else		
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else					
			credit_i(SOUTH) when tab_in(WEST)="011" and data_av(WEST)='1' else
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_av(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else
			data_in(WEST)  when tab_out(SOUTH)="001" and free(SOUTH)='0' else			
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmNLM;
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------------------
architecture AlgorithmNFM of Hermes_crossbar_TC is

begin
	tx(NORTH) <= '0';
	data_out(NORTH) <= (others=>'0');
	data_ack(NORTH) <= '0';
----------------------------------------------------------------------------------
-- PORTA LOCAL
----------------------------------------------------------------------------------
	tx(LOCAL) <= data_av(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_av(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_av(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			'0';

	data_out(LOCAL) <= data_in(EAST) when tab_out(LOCAL)="000" and free(LOCAL)='0' else
			data_in(WEST)  when tab_out(LOCAL)="001" and free(LOCAL)='0' else			
			data_in(SOUTH) when tab_out(LOCAL)="011" and free(LOCAL)='0' else
			(others=>'0');

	data_ack(LOCAL) <= credit_i(EAST) when tab_in(LOCAL)="000" and data_av(LOCAL)='1' else
			credit_i(WEST)  when tab_in(LOCAL)="001" and data_av(LOCAL)='1' else			
			credit_i(SOUTH) when tab_in(LOCAL)="011" and data_av(LOCAL)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA EAST
----------------------------------------------------------------------------------
	tx(EAST) <= data_av(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_av(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_av(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			'0';

	data_out(EAST) <= data_in(WEST) when tab_out(EAST)="001" and free(EAST)='0' else			
			data_in(SOUTH) when tab_out(EAST)="011" and free(EAST)='0' else
			data_in(LOCAL) when tab_out(EAST)="100" and free(EAST)='0' else
			(others=>'0');

	data_ack(EAST) <= credit_i(WEST) when tab_in(EAST)="001" and data_av(EAST)='1' else			
			credit_i(SOUTH) when tab_in(EAST)="011" and data_av(EAST)='1' else
			credit_i(LOCAL) when tab_in(EAST)="100" and data_av(EAST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA WEST
----------------------------------------------------------------------------------
	tx(WEST) <= data_av(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_av(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			'0';

	data_out(WEST) <= data_in(EAST) when tab_out(WEST)="000" and free(WEST)='0' else			
			data_in(LOCAL) when tab_out(WEST)="100" and free(WEST)='0' else
			(others=>'0');

	data_ack(WEST) <= credit_i(EAST) when tab_in(WEST)="000" and data_av(WEST)='1' else			
			credit_i(LOCAL) when tab_in(WEST)="100" and data_av(WEST)='1' else
			'0';
----------------------------------------------------------------------------------
-- PORTA SOUTH
----------------------------------------------------------------------------------
	tx(SOUTH) <= data_av(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else			
			data_av(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			'0';

	data_out(SOUTH) <= data_in(EAST) when tab_out(SOUTH)="000" and free(SOUTH)='0' else			
			data_in(LOCAL) when tab_out(SOUTH)="100" and free(SOUTH)='0' else
			(others=>'0');

	data_ack(SOUTH) <= credit_i(EAST) when tab_in(SOUTH)="000" and data_av(SOUTH)='1' else			
			credit_i(LOCAL) when tab_in(SOUTH)="100" and data_av(SOUTH)='1' else
			'0';

end AlgorithmNFM;
