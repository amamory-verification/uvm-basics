package hermes_pkg_hdl;

   //`include "src/spi_typedefs_hdl.svh"

endpackage
