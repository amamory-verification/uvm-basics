class hermes_agent_cfg extends uvm_object;
`uvm_object_utils(hermes_agent_cfg)



endclass : hermes_agent_cfg
